`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12.08.2023 18:42:16
// Design Name: 
// Module Name: Keccakf
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



module Keccakf(string1 ,string2);
input [1599:0]string1;
output [1599:0] string2;
wire [63:0]a00,a01,a02,a03,a04;
wire [63:0]a10,a11,a12,a13,a14;
wire [63:0]a20,a21,a22,a23,a24;
wire [63:0]a30,a31,a32,a33,a34;
wire [63:0]a40,a41,a42,a43,a44;

wire [63:0]c00[23:0],c01[23:0],c02[23:0],c03[23:0],c04[23:0];
wire [63:0]c10[23:0],c11[23:0],c12[23:0],c13[23:0],c14[23:0];
wire [63:0]c20[23:0],c21[23:0],c22[23:0],c23[23:0],c24[23:0];
wire [63:0]c30[23:0],c31[23:0],c32[23:0],c33[23:0],c34[23:0];
wire [63:0]c40[23:0],c41[23:0],c42[23:0],c43[23:0],c44[23:0];

assign c00[0]=a00,c01[0]=a01,c02[0]=a02,c03[0]=a03,c04[0]=a04;
assign c10[0]=a10,c11[0]=a11,c12[0]=a12,c13[0]=a13,c14[0]=a14;
assign c20[0]=a20,c21[0]=a21,c22[0]=a22,c23[0]=a23,c24[0]=a24;
assign c30[0]=a30,c31[0]=a31,c32[0]=a32,c33[0]=a33,c34[0]=a34;
assign c40[0]=a40,c41[0]=a41,c42[0]=a42,c43[0]=a43,c44[0]=a44;

wire [63:0]d00,d01,d02,d03,d04;
wire [63:0]d10,d11,d12,d13,d14;
wire [63:0]d20,d21,d22,d23,d24;
wire [63:0]d30,d31,d32,d33,d34;
wire [63:0]d40,d41,d42,d43,d44;

stringtostate S1 (string1,a00,a01,a02,a03,a04,a10,a11,a12,a13,a14,a20,a21,a22,a23,a24,a30,a31,a32,a33,a34,a40,a41,a42,a43,a44);
genvar i;

for(i=0;i<23;i=i+1)
begin
round A1(c00[i],c01[i],c02[i],c03[i],c04[i],c10[i],c11[i],c12[i],c13[i],c14[i],c20[i],c21[i],c22[i],c23[i],c24[i],c30[i],c31[i],c32[i],c33[i],c34[i],c40[i],c41[i],c42[i],c43[i],c44[i],
c00[i+1],c01[i+1],c02[i+1],c03[i+1],c04[i+1],c10[i+1],c11[i+1],c12[i+1],c13[i+1],c14[i+1],c20[i+1],c21[i+1],c22[i+1],c23[i+1],c24[i+1],c30[i+1],c31[i+1],c32[i+1],c33[i+1],c34[i+1],c40[i+1],c41[i+1],c42[i+1],c43[i+1],c44[i+1],i);

end

round A2(c00[23],c01[23],c02[23],c03[23],c04[23],c10[23],c11[23],c12[23],c13[23],c14[23],c20[23],c21[23],c22[23],c23[23],c24[23],c30[23],c31[23],c32[23],c33[23],c34[23],c40[23],c41[23],c42[23],c43[23],c44[23],
d00,d01,d02,d03,d04,d10,d11,d12,d13,d14,d20,d21,d22,d23,d24,d30,d31,d32,d33,d34,d40,d41,d42,d43,d44,23);

statetostring O1 (d00,d01,d02,d03,d04,d10,d11,d12,d13,d14,d20,d21,d22,d23,d24,d30,d31,d32,d33,d34,d40,d41,d42,d43,d44,string2);
endmodule
