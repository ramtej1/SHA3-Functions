`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 14.08.2023 12:37:51
// Design Name: 
// Module Name: thota
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module thota(a00,a01,a02,a03,a04,a10,a11,a12,a13,a14,a20,a21,a22,a23,a24,a30,a31,a32,a33,a34,a40,a41,a42,a43,a44,
b00,b01,b02,b03,b04,b10,b11,b12,b13,b14,b20,b21,b22,b23,b24,b30,b31,b32,b33,b34,b40,b41,b42,b43,b44
,ir
    );
    
input [63:0]a00,a01,a02,a03,a04;
input [63:0]a10,a11,a12,a13,a14;
input [63:0]a20,a21,a22,a23,a24;
input [63:0]a30,a31,a32,a33,a34;
input [63:0]a40,a41,a42,a43,a44;
input [31:0]ir;
  
output [63:0]b00,b01,b02,b03,b04;
output [63:0]b10,b11,b12,b13,b14;
output [63:0]b20,b21,b22,b23,b24;
output [63:0]b30,b31,b32,b33,b34;
output [63:0]b40,b41,b42,b43,b44;
genvar i;
wire [63:0] rc;
assign rc= ir==0?64'h0000000000000001:ir==1?64'h0000000000008082:ir==2?64'h800000000000808a:
ir==3?64'h8000000080008000:ir==4?64'h000000000000808b:ir==5?64'h0000000080000001:
ir==6?64'h8000000080008081:ir==7?64'h8000000000008009:ir==8?64'h000000000000008a:ir==9?64'h0000000000000088
:ir==10?64'h0000000080008009:ir==11?64'h000000008000000a:ir==12?64'h000000008000808b:
ir==13?64'h800000000000008b:ir==14?64'h8000000000008089:ir==15?64'h8000000000008003:
ir==16?64'h8000000000008002:ir==17?64'h8000000000000080:ir==18?64'h000000000000800a:
ir==19?64'h800000008000000a:ir==20?64'h8000000080008081:ir==21?64'h8000000000008080:
ir==22?64'h0000000080000001:ir==23?64'h8000000080008008:0;


assign b00 = a00^rc,b01 = a01,b02 = a02,b03 = a03,b04 = a04;
assign b10 = a10,b11 = a11,b12 = a12,b13 = a13,b14 = a14;
assign b20 = a20,b21 = a21,b22 = a22,b23 = a23,b24 = a24;
assign b30 = a30,b31 = a31,b32 = a32,b33 = a33,b34 = a34;
assign b40 = a40,b41 = a41,b42 = a42,b43 = a43,b44 = a44;
endmodule
